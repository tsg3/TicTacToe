module matrix_memory(input [3:0] m_cell, [1:0] player, aceptar, clk, rst, output [4:0] next_play);